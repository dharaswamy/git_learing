
/*

File Name : apb_scoreboard.sv
Purpose   : It is a reference model and it will check the Actual vlaues with expected values ang give whether the test is passed or failed . 

*/ 

class apb_scoreboard extends uvm_scrorboard;

  //uvm Factory registration
  uvm_component_utils(apb_scoreboard) 

  
endclass:apb_scoreboard 

