
/*

File Name : apb_subscriber.sv
Purpose   : It measure functional coverage of apb protocol .

*/

class apb_subscriber extends uvm_subscriber#(apb_sequence_item);

  //Factory Registration
   uvm_component_utils(apb_subscriber) 


endclass:apb_subscriber


